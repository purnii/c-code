module ha(sum,car,a,b);
  input a,b;
  output sum,car;
  wire a;
  wire b;
  reg sum;
  reg car;
  ha(sum,car,a,b);
endmodule
  
