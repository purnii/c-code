module fa(sum,car,a,b);
  input a,b;
  output sum,car;
  wire a;
  wire b;
  wire sum;
  wire car;
  ha(sum,car,a,b);
endmodule

