module three_to_8_decoder(z,x0,x1,x2);
  input x0,x1,x2;
  output [7:0]z;
  wire p0,p1,p2;
  not (p0,x0);
  not (p1,x1);
  not (p2,x2);
  and (z[0],p2,p1,p0);
  and (z[1],p2,p1,x0);
  and (z[2],p2,x1,p0);
  and (z[3],p2,x1,x0);
  and (z[4],x2,p1,p0);
  and (z[5],x2,p1,x0);
  and (z[6],x2,x1,p0);
  and (z[7],x2,x1,x0);
endmodule
